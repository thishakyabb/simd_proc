`ifndef PARAMS_SVH
`define PARAMS_SVH

parameter OP_SEL_WIDTH = 2;
parameter OPCODE_WIDTH = 3;

`endif